module unidad_control();

endmodule 