module registro_MEM_WB();

endmodule
