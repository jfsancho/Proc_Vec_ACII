module registro_EXE_MEM();

endmodule
