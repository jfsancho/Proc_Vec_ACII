// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: mux_8x10.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 16.1.0 Build 196 10/24/2016 SJ Lite Edition
// ************************************************************


//Copyright (C) 2016  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Intel and sold by Intel or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module mux_8x10 (
	data0x,
	data1x,
	data2x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	sel,
	result);

	input	[9:0]  data0x;
	input	[9:0]  data1x;
	input	[9:0]  data2x;
	input	[9:0]  data3x;
	input	[9:0]  data4x;
	input	[9:0]  data5x;
	input	[9:0]  data6x;
	input	[9:0]  data7x;
	input	[2:0]  sel;
	output	[9:0]  result;

	wire [9:0] sub_wire9;
	wire [9:0] sub_wire8 = data7x[9:0];
	wire [9:0] sub_wire7 = data6x[9:0];
	wire [9:0] sub_wire6 = data5x[9:0];
	wire [9:0] sub_wire5 = data4x[9:0];
	wire [9:0] sub_wire4 = data3x[9:0];
	wire [9:0] sub_wire3 = data2x[9:0];
	wire [9:0] sub_wire2 = data1x[9:0];
	wire [9:0] sub_wire0 = data0x[9:0];
	wire [79:0] sub_wire1 = {sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire2, sub_wire0};
	wire [9:0] result = sub_wire9[9:0];

	lpm_mux	LPM_MUX_component (
				.data (sub_wire1),
				.sel (sel),
				.result (sub_wire9)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_size = 8,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = 10,
		LPM_MUX_component.lpm_widths = 3;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone V"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "8"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "10"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "3"
// Retrieval info: USED_PORT: data0x 0 0 10 0 INPUT NODEFVAL "data0x[9..0]"
// Retrieval info: USED_PORT: data1x 0 0 10 0 INPUT NODEFVAL "data1x[9..0]"
// Retrieval info: USED_PORT: data2x 0 0 10 0 INPUT NODEFVAL "data2x[9..0]"
// Retrieval info: USED_PORT: data3x 0 0 10 0 INPUT NODEFVAL "data3x[9..0]"
// Retrieval info: USED_PORT: data4x 0 0 10 0 INPUT NODEFVAL "data4x[9..0]"
// Retrieval info: USED_PORT: data5x 0 0 10 0 INPUT NODEFVAL "data5x[9..0]"
// Retrieval info: USED_PORT: data6x 0 0 10 0 INPUT NODEFVAL "data6x[9..0]"
// Retrieval info: USED_PORT: data7x 0 0 10 0 INPUT NODEFVAL "data7x[9..0]"
// Retrieval info: USED_PORT: result 0 0 10 0 OUTPUT NODEFVAL "result[9..0]"
// Retrieval info: USED_PORT: sel 0 0 3 0 INPUT NODEFVAL "sel[2..0]"
// Retrieval info: CONNECT: @data 0 0 10 0 data0x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 10 data1x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 20 data2x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 30 data3x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 40 data4x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 50 data5x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 60 data6x 0 0 10 0
// Retrieval info: CONNECT: @data 0 0 10 70 data7x 0 0 10 0
// Retrieval info: CONNECT: @sel 0 0 3 0 sel 0 0 3 0
// Retrieval info: CONNECT: result 0 0 10 0 @result 0 0 10 0
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL mux_8x10_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
